`timescale 1ns/1ps

module tb_shift_add_multiplier;

    // Sinais
    logic clk;
    logic rst;
    logic [7:0] multiplicand;
    logic [7:0] multiplier;
    logic [15:0] result;
    logic end_op;

    // DUT
    shift_add_multiplier uut (
        .clk(clk), .rst(rst), .multiplicand(multiplicand), .multiplier(multiplier),
        .result(result), .end_op(end_op)
    );

    // Clock 10 ns
    initial clk = 0;
    always #5 clk = ~clk;

    // Vetores de teste
    logic [7:0] test_a [0:5];
    logic [7:0] test_b [0:5];

    integer i;
    integer cycles;
    integer timeout;
    logic [15:0] expected;

    initial begin
    // grava o VCD na pasta sim do projeto mesmo quando a simula                                   
    $dumpfile("../sim/shift_add_multiplier.vcd");
        $dumpvars(0, tb_shift_add_multiplier);

        // Vetores
        test_a[0] = 8'd3;   test_b[0] = 8'd5;
        test_a[1] = 8'd10;  test_b[1] = 8'd12;
        test_a[2] = 8'd127; test_b[2] = 8'd201;
        test_a[3] = 8'd255; test_b[3] = 8'd255;
        test_a[4] = 8'd0;   test_b[4] = 8'd123;
        test_a[5] = 8'd13;  test_b[5] = 8'd11;

    // Loop de testes
        for (i = 0; i < 6; i = i + 1) begin
            multiplicand = test_a[i];
            multiplier   = test_b[i];

            // Reset do DUT
            rst = 1;
            @(posedge clk);
            @(posedge clk);
            rst = 0;

            // Espera fim ou timeout
            cycles = 0;
            timeout = 200;
            while (!end_op && cycles < timeout) begin
                    @(posedge clk);
                    cycles = cycles + 1;
                    // Debug interno
                    $display(" ciclo=%0d estado=%0d cnt=%0d A=0x%0h B=0x%0h Q=0x%0h | soma=0x%0h c_out=%b",
                        cycles, uut.state, uut.iter_cnt.data_out, uut.A_out, uut.B_out, uut.Q_out, uut.sum, uut.c_out);
            end

            // Resultado esperado
            expected = multiplicand * multiplier;

            $display("--------------------------------------------------");
            $display("Teste %0d: %0d x %0d", i, multiplicand, multiplier);
            $display("Ciclos aguardados: %0d, fim=%0b", cycles, end_op);
            $display("Resultado DUT = %0d (0x%0h), Esperado = %0d (0x%0h)", result, result, expected, expected);
            if (result === expected) $display("OK"); else $display("FALHOU");

            // Espaço entre testes
            repeat (4) @(posedge clk);
        end

    $display("Todos os testes concluidos.");
        #20 $finish;
    end

endmodule
